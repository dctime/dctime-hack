module hack( input in, output out );
	assign out = ~in;
endmodule