module And (
    input in_a,
    input in_b,
    output out_a
);

assign out_a = in_a & in_b;
    
endmodule